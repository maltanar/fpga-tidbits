module GenericSDAccelWrapperTop(input clk, input reset,
    output s_axi_control_AWREADY,
    input  s_axi_control_AWVALID,
    input [63:0] s_axi_control_AWADDR,
    input [2:0] s_axi_control_AWPROT,
    output s_axi_control_WREADY,
    input  s_axi_control_WVALID,
    input [31:0] s_axi_control_WDATA,
    input [3:0] s_axi_control_WSTRB,
    input  s_axi_control_BREADY,
    output s_axi_control_BVALID,
    output[1:0] s_axi_control_BRESP,
    output s_axi_control_ARREADY,
    input  s_axi_control_ARVALID,
    input [63:0] s_axi_control_ARADDR,
    input [2:0] s_axi_control_ARPROT,
    input  s_axi_control_RREADY,
    output s_axi_control_RVALID,
    output[31:0] s_axi_control_RDATA,
    output[1:0] s_axi_control_RRESP,
    input  mem0_AWREADY,
    output mem0_AWVALID,
    output[63:0] mem0_AWADDR,
    output[2:0] mem0_AWSIZE,
    output[7:0] mem0_AWLEN,
    output[1:0] mem0_AWBURST,
    output[5:0] mem0_AWID,
    output mem0_AWLOCK,
    output[3:0] mem0_AWCACHE,
    output[2:0] mem0_AWPROT,
    output[3:0] mem0_AWQOS,
    input  mem0_WREADY,
    output mem0_WVALID,
    output[511:0] mem0_WDATA,
    output[63:0] mem0_WSTRB,
    output mem0_WLAST,
    output mem0_BREADY,
    input  mem0_BVALID,
    input [5:0] mem0_BID,
    input [1:0] mem0_BRESP,
    input  mem0_ARREADY,
    output mem0_ARVALID,
    output[63:0] mem0_ARADDR,
    output[2:0] mem0_ARSIZE,
    output[7:0] mem0_ARLEN,
    output[1:0] mem0_ARBURST,
    output[5:0] mem0_ARID,
    output mem0_ARLOCK,
    output[3:0] mem0_ARCACHE,
    output[2:0] mem0_ARPROT,
    output[3:0] mem0_ARQOS,
    output mem0_RREADY,
    input  mem0_RVALID,
    input [511:0] mem0_RDATA,
    input [5:0] mem0_RID,
    input  mem0_RLAST,
    input [1:0] mem0_RRESP
);
  GenericSDAccelWrapper GenericSDAccelWrapper(.clk(ap_clk), .reset(!ap_rst_n),
  	.csr_AWREADY(s_axi_control_AWREADY),
		.csr_AWVALID(s_axi_control_AWVALID),
		.csr_AWADDR(s_axi_control_AWADDR),
		.csr_AWPROT(s_axi_control_AWPROT),
		.csr_WREADY(s_axi_control_WREADY),
		.csr_WVALID(s_axi_control_WVALID),
		.csr_WDATA(s_axi_control_WDATA),
		.csr_WSTRB(s_axi_control_WSTRB),
		.csr_BREADY(s_axi_control_BREADY),
		.csr_BVALID(s_axi_control_BVALID),
		.csr_BRESP(s_axi_control_BRESP),
		.csr_ARREADY(s_axi_control_ARREADY),
		.csr_ARVALID(s_axi_control_ARVALID),
		.csr_ARADDR(s_axi_control_ARADDR),
		.csr_ARPROT(s_axi_control_ARPROT),
		.csr_RREADY(s_axi_control_RREADY),
		.csr_RVALID(s_axi_control_RVALID),
		.csr_RDATA(s_axi_control_RDATA),
		.csr_RRESP(s_axi_control_RRESP),
		.mem0_AWREADY(mem0_AWREADY),
		.mem0_AWVALID(mem0_AWVALID),
		.mem0_AWADDR(mem0_AWADDR),
		.mem0_AWSIZE(mem0_AWSIZE),
		.mem0_AWLEN(mem0_AWLEN),
		.mem0_AWBURST(mem0_AWBURST),
		.mem0_AWID(mem0_AWID),
		.mem0_AWLOCK(mem0_AWLOCK),
		.mem0_AWCACHE(mem0_AWCACHE),
		.mem0_AWPROT(mem0_AWPROT),
		.mem0_AWQOS(mem0_AWQOS),
		.mem0_WREADY(mem0_WREADY),
		.mem0_WVALID(mem0_WVALID),
		.mem0_WDATA(mem0_WDATA),
		.mem0_WSTRB(mem0_WSTRB),
		.mem0_WLAST(mem0_WLAST),
		.mem0_BREADY(mem0_BREADY),
		.mem0_BVALID(mem0_BVALID),
		.mem0_BID(mem0_BID),
		.mem0_BRESP(mem0_BRESP),
		.mem0_ARREADY(mem0_ARREADY),
		.mem0_ARVALID(mem0_ARVALID),
		.mem0_ARADDR(mem0_ARADDR),
		.mem0_ARSIZE(mem0_ARSIZE),
		.mem0_ARLEN(mem0_ARLEN),
		.mem0_ARBURST(mem0_ARBURST),
		.mem0_ARID(mem0_ARID),
		.mem0_ARLOCK(mem0_ARLOCK),
		.mem0_ARCACHE(mem0_ARCACHE),
		.mem0_ARPROT(mem0_ARPROT),
		.mem0_ARQOS(mem0_ARQOS),
		.mem0_RREADY(mem0_RREADY),
		.mem0_RVALID(mem0_RVALID),
		.mem0_RDATA(mem0_RDATA),
		.mem0_RID(mem0_RID),
		.mem0_RLAST(mem0_RLAST),
		.mem0_RRESP(mem0_RRESP)
  );
endmodule
