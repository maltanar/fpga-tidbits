module ZedBoardWrapper(input clk, input reset,
    output csr_AWREADY,
    input  csr_AWVALID,
    input [31:0] csr_AWADDR,
    input [2:0] csr_AWPROT,
    output csr_WREADY,
    input  csr_WVALID,
    input [31:0] csr_WDATA,
    input [3:0] csr_WSTRB,
    input  csr_BREADY,
    output csr_BVALID,
    output[1:0] csr_BRESP,
    output csr_ARREADY,
    input  csr_ARVALID,
    input [31:0] csr_ARADDR,
    input [2:0] csr_ARPROT,
    input  csr_RREADY,
    output csr_RVALID,
    output[31:0] csr_RDATA,
    output[1:0] csr_RRESP,
    input  mem3_AWREADY,
    output mem3_AWVALID,
    output[31:0] mem3_AWADDR,
    output[2:0] mem3_AWSIZE,
    output[7:0] mem3_AWLEN,
    output[1:0] mem3_AWBURST,
    output[5:0] mem3_AWID,
    output mem3_AWLOCK,
    output[3:0] mem3_AWCACHE,
    output[2:0] mem3_AWPROT,
    output[3:0] mem3_AWQOS,
    input  mem3_WREADY,
    output mem3_WVALID,
    output[63:0] mem3_WDATA,
    output[7:0] mem3_WSTRB,
    output mem3_WLAST,
    output mem3_BREADY,
    input  mem3_BVALID,
    input [5:0] mem3_BID,
    input [1:0] mem3_BRESP,
    input  mem3_ARREADY,
    output mem3_ARVALID,
    output[31:0] mem3_ARADDR,
    output[2:0] mem3_ARSIZE,
    output[7:0] mem3_ARLEN,
    output[1:0] mem3_ARBURST,
    output[5:0] mem3_ARID,
    output mem3_ARLOCK,
    output[3:0] mem3_ARCACHE,
    output[2:0] mem3_ARPROT,
    output[3:0] mem3_ARQOS,
    output mem3_RREADY,
    input  mem3_RVALID,
    input [63:0] mem3_RDATA,
    input [5:0] mem3_RID,
    input  mem3_RLAST,
    input [1:0] mem3_RRESP,
    input  mem2_AWREADY,
    output mem2_AWVALID,
    output[31:0] mem2_AWADDR,
    output[2:0] mem2_AWSIZE,
    output[7:0] mem2_AWLEN,
    output[1:0] mem2_AWBURST,
    output[5:0] mem2_AWID,
    output mem2_AWLOCK,
    output[3:0] mem2_AWCACHE,
    output[2:0] mem2_AWPROT,
    output[3:0] mem2_AWQOS,
    input  mem2_WREADY,
    output mem2_WVALID,
    output[63:0] mem2_WDATA,
    output[7:0] mem2_WSTRB,
    output mem2_WLAST,
    output mem2_BREADY,
    input  mem2_BVALID,
    input [5:0] mem2_BID,
    input [1:0] mem2_BRESP,
    input  mem2_ARREADY,
    output mem2_ARVALID,
    output[31:0] mem2_ARADDR,
    output[2:0] mem2_ARSIZE,
    output[7:0] mem2_ARLEN,
    output[1:0] mem2_ARBURST,
    output[5:0] mem2_ARID,
    output mem2_ARLOCK,
    output[3:0] mem2_ARCACHE,
    output[2:0] mem2_ARPROT,
    output[3:0] mem2_ARQOS,
    output mem2_RREADY,
    input  mem2_RVALID,
    input [63:0] mem2_RDATA,
    input [5:0] mem2_RID,
    input  mem2_RLAST,
    input [1:0] mem2_RRESP,
    input  mem1_AWREADY,
    output mem1_AWVALID,
    output[31:0] mem1_AWADDR,
    output[2:0] mem1_AWSIZE,
    output[7:0] mem1_AWLEN,
    output[1:0] mem1_AWBURST,
    output[5:0] mem1_AWID,
    output mem1_AWLOCK,
    output[3:0] mem1_AWCACHE,
    output[2:0] mem1_AWPROT,
    output[3:0] mem1_AWQOS,
    input  mem1_WREADY,
    output mem1_WVALID,
    output[63:0] mem1_WDATA,
    output[7:0] mem1_WSTRB,
    output mem1_WLAST,
    output mem1_BREADY,
    input  mem1_BVALID,
    input [5:0] mem1_BID,
    input [1:0] mem1_BRESP,
    input  mem1_ARREADY,
    output mem1_ARVALID,
    output[31:0] mem1_ARADDR,
    output[2:0] mem1_ARSIZE,
    output[7:0] mem1_ARLEN,
    output[1:0] mem1_ARBURST,
    output[5:0] mem1_ARID,
    output mem1_ARLOCK,
    output[3:0] mem1_ARCACHE,
    output[2:0] mem1_ARPROT,
    output[3:0] mem1_ARQOS,
    output mem1_RREADY,
    input  mem1_RVALID,
    input [63:0] mem1_RDATA,
    input [5:0] mem1_RID,
    input  mem1_RLAST,
    input [1:0] mem1_RRESP,
    input  mem0_AWREADY,
    output mem0_AWVALID,
    output[31:0] mem0_AWADDR,
    output[2:0] mem0_AWSIZE,
    output[7:0] mem0_AWLEN,
    output[1:0] mem0_AWBURST,
    output[5:0] mem0_AWID,
    output mem0_AWLOCK,
    output[3:0] mem0_AWCACHE,
    output[2:0] mem0_AWPROT,
    output[3:0] mem0_AWQOS,
    input  mem0_WREADY,
    output mem0_WVALID,
    output[63:0] mem0_WDATA,
    output[7:0] mem0_WSTRB,
    output mem0_WLAST,
    output mem0_BREADY,
    input  mem0_BVALID,
    input [5:0] mem0_BID,
    input [1:0] mem0_BRESP,
    input  mem0_ARREADY,
    output mem0_ARVALID,
    output[31:0] mem0_ARADDR,
    output[2:0] mem0_ARSIZE,
    output[7:0] mem0_ARLEN,
    output[1:0] mem0_ARBURST,
    output[5:0] mem0_ARID,
    output mem0_ARLOCK,
    output[3:0] mem0_ARCACHE,
    output[2:0] mem0_ARPROT,
    output[3:0] mem0_ARQOS,
    output mem0_RREADY,
    input  mem0_RVALID,
    input [63:0] mem0_RDATA,
    input [5:0] mem0_RID,
    input  mem0_RLAST,
    input [1:0] mem0_RRESP
);


endmodule