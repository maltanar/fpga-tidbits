module GenericSDAccelWrapperTop(input ap_clk, input ap_rst_n,
    output s_axi_control_AWREADY,
    input  s_axi_control_AWVALID,
    input [63:0] s_axi_control_AWADDR,
    input [2:0] s_axi_control_AWPROT,
    output s_axi_control_WREADY,
    input  s_axi_control_WVALID,
    input [31:0] s_axi_control_WDATA,
    input [3:0] s_axi_control_WSTRB,
    input  s_axi_control_BREADY,
    output s_axi_control_BVALID,
    output[1:0] s_axi_control_BRESP,
    output s_axi_control_ARREADY,
    input  s_axi_control_ARVALID,
    input [63:0] s_axi_control_ARADDR,
    input [2:0] s_axi_control_ARPROT,
    input  s_axi_control_RREADY,
    output s_axi_control_RVALID,
    output[31:0] s_axi_control_RDATA,
    output[1:0] s_axi_control_RRESP,
    input  m_axi_gmem_AWREADY,
    output m_axi_gmem_AWVALID,
    output[63:0] m_axi_gmem_AWADDR,
    output[2:0] m_axi_gmem_AWSIZE,
    output[7:0] m_axi_gmem_AWLEN,
    output[1:0] m_axi_gmem_AWBURST,
    output[0:0] m_axi_gmem_AWID,
    output m_axi_gmem_AWLOCK,
    output[3:0] m_axi_gmem_AWCACHE,
    output[2:0] m_axi_gmem_AWPROT,
    output[3:0] m_axi_gmem_AWQOS,
    input  m_axi_gmem_WREADY,
    output m_axi_gmem_WVALID,
    output[63:0] m_axi_gmem_WDATA,
    output[63:0] m_axi_gmem_WSTRB,
    output m_axi_gmem_WLAST,
    output m_axi_gmem_BREADY,
    input  m_axi_gmem_BVALID,
    input [0:0] m_axi_gmem_BID,
    input [1:0] m_axi_gmem_BRESP,
    input  m_axi_gmem_ARREADY,
    output m_axi_gmem_ARVALID,
    output[63:0] m_axi_gmem_ARADDR,
    output[2:0] m_axi_gmem_ARSIZE,
    output[7:0] m_axi_gmem_ARLEN,
    output[1:0] m_axi_gmem_ARBURST,
    output[0:0] m_axi_gmem_ARID,
    output m_axi_gmem_ARLOCK,
    output[3:0] m_axi_gmem_ARCACHE,
    output[2:0] m_axi_gmem_ARPROT,
    output[3:0] m_axi_gmem_ARQOS,
    output m_axi_gmem_RREADY,
    input  m_axi_gmem_RVALID,
    input [63:0] m_axi_gmem_RDATA,
    input [0:0] m_axi_gmem_RID,
    input  m_axi_gmem_RLAST,
    input [1:0] m_axi_gmem_RRESP
);
  GenericSDAccelWrapper GenericSDAccelWrapper(.clk(ap_clk), .reset(!ap_rst_n),
  	.csr_AWREADY(s_axi_control_AWREADY),
		.csr_AWVALID(s_axi_control_AWVALID),
		.csr_AWADDR(s_axi_control_AWADDR),
		.csr_AWPROT(s_axi_control_AWPROT),
		.csr_WREADY(s_axi_control_WREADY),
		.csr_WVALID(s_axi_control_WVALID),
		.csr_WDATA(s_axi_control_WDATA),
		.csr_WSTRB(s_axi_control_WSTRB),
		.csr_BREADY(s_axi_control_BREADY),
		.csr_BVALID(s_axi_control_BVALID),
		.csr_BRESP(s_axi_control_BRESP),
		.csr_ARREADY(s_axi_control_ARREADY),
		.csr_ARVALID(s_axi_control_ARVALID),
		.csr_ARADDR(s_axi_control_ARADDR),
		.csr_ARPROT(s_axi_control_ARPROT),
		.csr_RREADY(s_axi_control_RREADY),
		.csr_RVALID(s_axi_control_RVALID),
		.csr_RDATA(s_axi_control_RDATA),
		.csr_RRESP(s_axi_control_RRESP),
		.mem0_AWREADY(m_axi_gmem_AWREADY),
		.mem0_AWVALID(m_axi_gmem_AWVALID),
		.mem0_AWADDR(m_axi_gmem_AWADDR),
		.mem0_AWSIZE(m_axi_gmem_AWSIZE),
		.mem0_AWLEN(m_axi_gmem_AWLEN),
		.mem0_AWBURST(m_axi_gmem_AWBURST),
		.mem0_AWID(m_axi_gmem_AWID),
		.mem0_AWLOCK(m_axi_gmem_AWLOCK),
		.mem0_AWCACHE(m_axi_gmem_AWCACHE),
		.mem0_AWPROT(m_axi_gmem_AWPROT),
		.mem0_AWQOS(m_axi_gmem_AWQOS),
		.mem0_WREADY(m_axi_gmem_WREADY),
		.mem0_WVALID(m_axi_gmem_WVALID),
		.mem0_WDATA(m_axi_gmem_WDATA),
		.mem0_WSTRB(m_axi_gmem_WSTRB),
		.mem0_WLAST(m_axi_gmem_WLAST),
		.mem0_BREADY(m_axi_gmem_BREADY),
		.mem0_BVALID(m_axi_gmem_BVALID),
		.mem0_BID(m_axi_gmem_BID),
		.mem0_BRESP(m_axi_gmem_BRESP),
		.mem0_ARREADY(m_axi_gmem_ARREADY),
		.mem0_ARVALID(m_axi_gmem_ARVALID),
		.mem0_ARADDR(m_axi_gmem_ARADDR),
		.mem0_ARSIZE(m_axi_gmem_ARSIZE),
		.mem0_ARLEN(m_axi_gmem_ARLEN),
		.mem0_ARBURST(m_axi_gmem_ARBURST),
		.mem0_ARID(m_axi_gmem_ARID),
		.mem0_ARLOCK(m_axi_gmem_ARLOCK),
		.mem0_ARCACHE(m_axi_gmem_ARCACHE),
		.mem0_ARPROT(m_axi_gmem_ARPROT),
		.mem0_ARQOS(m_axi_gmem_ARQOS),
		.mem0_RREADY(m_axi_gmem_RREADY),
		.mem0_RVALID(m_axi_gmem_RVALID),
		.mem0_RDATA(m_axi_gmem_RDATA),
		.mem0_RID(m_axi_gmem_RID),
		.mem0_RLAST(m_axi_gmem_RLAST),
		.mem0_RRESP(m_axi_gmem_RRESP)
  );
endmodule
